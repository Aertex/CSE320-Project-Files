This is a test to see if git recognizes systemverilog aka .sv files