`timescale 1ns / 1ps

//just holds container, 
module TopModule(
input logic switch0,
input logic switch1,
input logic reset,
input logic play,
input logic record,

input logic microphone,
output logic audio_out,

output logic a0,
output logic a1,
output logic [6:0]cathode

    );




endmodule