`timescale 1ns / 1ps
//reads input from microphone, stores it into memory
//needs to read a line of 0/1 and creates a 16 bit word
//outputs done signal every 16 clock cycles
//needs to convert a 100mhz clock signal to 1mhz signal internally
module Deserializer(

    );
endmodule
